module NegativeFlag (input logic LB,
					  output logic Res);
										
	assign Res = LB;

endmodule 