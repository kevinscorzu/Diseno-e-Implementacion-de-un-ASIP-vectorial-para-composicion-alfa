//module PipelineDecode()

//endmodule 